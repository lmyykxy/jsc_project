 //`define sim
`define project